CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 120 30 70 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
37
13 Logic Switch~
5 364 640 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8585 0 0
2
5.90072e-315 0
0
13 Logic Switch~
5 310 638 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8809 0 0
2
5.90072e-315 0
0
8 2-In OR~
219 85 615 0 3 22
0 5 23 17
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U1C
-5 20 16 28
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5993 0 0
2
5.90072e-315 0
0
9 Inverter~
13 180 615 0 2 22
0 17 21
0
0 0 624 0
5 74F04
-18 -19 17 -11
4 U19A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 10 0
1 U
8654 0 0
2
5.90072e-315 0
0
9 2-In AND~
219 237 606 0 3 22
0 6 21 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
7223 0 0
2
5.90072e-315 0
0
6 74LS47
187 1671 267 0 14 29
0 33 36 32 35 86 87 34 44 45
46 47 48 49 88
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
3 U17
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3641 0 0
2
5.90072e-315 5.37752e-315
0
9 CA 7-Seg~
184 1729 161 0 18 19
10 49 48 47 46 45 44 34 89 90
0 0 0 0 0 0 0 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3104 0 0
2
5.90072e-315 5.36716e-315
0
6 74LS93
109 1565 240 0 8 17
0 26 26 19 35 33 36 32 35
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
3 U16
-10 -36 11 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3296 0 0
2
5.90072e-315 5.3568e-315
0
6 74LS93
109 1310 249 0 8 17
0 20 20 26 30 31 28 29 30
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
3 U15
-10 -36 11 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
8534 0 0
2
5.90072e-315 5.34643e-315
0
9 CA 7-Seg~
184 1462 158 0 18 19
10 43 42 41 40 39 38 37 91 92
2 0 0 2 2 2 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
949 0 0
2
5.90072e-315 5.32571e-315
0
6 74LS47
187 1394 276 0 14 29
0 31 28 29 30 93 94 37 38 39
40 41 42 43 95
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
3 U14
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3371 0 0
2
5.90072e-315 5.30499e-315
0
9 2-In AND~
219 1511 338 0 3 22
0 32 33 26
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 U13C
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
7311 0 0
2
5.90072e-315 5.26354e-315
0
9 2-In AND~
219 1266 377 0 3 22
0 29 28 20
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 U13B
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3409 0 0
2
5.90072e-315 0
0
9 2-In AND~
219 703 385 0 3 22
0 10 11 18
0
0 0 624 90
5 74F08
-18 -24 17 -16
4 U13A
13 -5 41 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
3526 0 0
2
5.90072e-315 0
0
9 2-In AND~
219 979 378 0 3 22
0 13 14 12
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U5D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
4129 0 0
2
5.90072e-315 0
0
7 Pulser~
4 1452 443 0 10 12
0 27 96 19 97 0 0 5 5 5
8
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6278 0 0
2
45027.4 0
0
6 74LS47
187 890 283 0 14 29
0 50 11 10 9 98 99 52 53 54
55 56 57 58 100
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
3 U12
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3482 0 0
2
45027.4 1
0
9 CA 7-Seg~
184 961 173 0 18 19
10 58 57 56 55 54 53 52 101 102
0 0 0 0 2 2 0 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8323 0 0
2
45027.4 2
0
6 74LS93
109 760 256 0 8 17
0 18 18 12 9 50 11 10 9
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
3 U11
-10 -36 11 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3984 0 0
2
45027.4 3
0
6 74LS93
109 1050 238 0 8 17
0 12 12 20 15 16 14 13 15
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
3 U10
-10 -36 11 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
7622 0 0
2
45027.4 4
0
9 CA 7-Seg~
184 1242 167 0 18 19
10 64 63 62 61 60 59 51 103 104
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
816 0 0
2
45027.4 5
0
6 74LS47
187 1175 265 0 14 29
0 16 14 13 15 105 106 51 59 60
61 62 63 64 107
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4656 0 0
2
45027.4 6
0
9 2-In AND~
219 175 533 0 3 22
0 7 6 65
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
6356 0 0
2
5.90072e-315 5.30499e-315
0
14 Logic Display~
6 551 532 0 1 2
12 66
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7479 0 0
2
5.90072e-315 5.32571e-315
0
9 2-In AND~
219 239 558 0 3 22
0 65 5 25
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
5690 0 0
2
5.90072e-315 5.34643e-315
0
6 74112~
219 311 594 0 7 32
0 2 25 18 22 24 108 66
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 6 0
1 U
5617 0 0
2
5.90072e-315 5.3568e-315
0
8 2-In OR~
219 333 320 0 3 22
0 68 67 69
0
0 0 624 90
5 74F32
-18 -24 17 -16
3 U1B
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3903 0 0
2
45027.4 7
0
9 2-In AND~
219 350 470 0 3 22
0 3 4 6
0
0 0 624 180
5 74F08
-18 -24 17 -16
3 U7D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4452 0 0
2
45027.4 9
0
9 2-In AND~
219 279 390 0 3 22
0 23 6 68
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U7C
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6282 0 0
2
45027.4 10
0
6 74LS93
109 185 240 0 8 17
0 68 68 67 5 71 70 23 5
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U9
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
7187 0 0
2
45027.4 12
0
6 74LS47
187 262 267 0 14 29
0 71 70 23 5 109 110 72 73 74
75 76 77 78 111
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6866 0 0
2
45027.4 13
0
9 CA 7-Seg~
184 323 183 0 18 19
10 78 77 76 75 74 73 72 112 113
0 0 0 0 0 0 2 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7670 0 0
2
45027.4 14
0
9 2-In AND~
219 346 393 0 3 22
0 8 7 67
0
0 0 624 90
5 74F08
-18 -24 17 -16
3 U7A
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
951 0 0
2
45027.4 15
0
6 74LS47
187 524 283 0 14 29
0 8 4 7 3 114 115 79 80 81
82 83 84 85 116
0
0 0 4848 0
7 74LS247
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9536 0 0
2
45027.4 16
0
9 CA 7-Seg~
184 581 179 0 18 19
10 85 84 83 82 81 80 79 117 118
2 2 0 0 0 0 0 2 2
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5495 0 0
2
45027.4 17
0
6 74LS93
109 419 256 0 8 17
0 69 69 18 3 8 4 7 3
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
8152 0 0
2
45027.4 18
0
2 +V
167 1402 427 0 1 3
0 27
0
0 0 54256 0
2 5V
-7 -24 7 -16
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6223 0 0
2
45027.4 19
0
122
1 1 2 0 0 4224 0 1 26 0 0 3
365 627
365 531
311 531
0 1 3 0 0 4224 0 0 28 6 0 3
448 289
448 479
368 479
0 2 4 0 0 4224 0 0 28 9 0 3
475 256
475 461
368 461
0 1 5 0 0 12432 0 0 3 90 0 5
106 429
106 427
43 427
43 606
72 606
2 0 6 0 0 4096 0 23 0 0 33 2
151 542
82 542
4 0 3 0 0 0 0 36 0 0 7 5
381 274
370 274
370 289
460 289
460 274
4 8 3 0 0 0 0 34 36 0 0 2
492 274
451 274
0 2 7 0 0 4096 0 0 33 115 0 4
469 265
469 439
354 439
354 414
6 2 4 0 0 0 0 36 34 0 0 2
451 256
492 256
1 0 8 0 0 12416 0 33 0 0 11 4
336 414
336 419
483 419
483 247
5 1 8 0 0 0 0 36 34 0 0 2
451 247
492 247
4 0 9 0 0 12416 0 19 0 0 13 5
722 274
711 274
711 289
802 289
802 274
8 4 9 0 0 0 0 19 17 0 0 2
792 274
858 274
1 0 10 0 0 12416 0 14 0 0 73 4
693 406
693 415
827 415
827 265
2 0 11 0 0 12416 0 14 0 0 74 4
711 406
711 410
847 410
847 256
3 0 12 0 0 12416 0 19 0 0 18 4
722 265
708 265
708 339
978 339
2 1 12 0 0 0 0 20 20 0 0 2
1018 238
1018 229
3 1 12 0 0 0 0 15 20 0 0 3
978 354
978 229
1018 229
1 0 13 0 0 12416 0 15 0 0 23 4
969 399
969 409
1114 409
1114 247
2 0 14 0 0 12416 0 15 0 0 24 4
987 399
987 404
1126 404
1126 238
4 8 15 0 0 12416 0 20 20 0 0 6
1012 256
1009 256
1009 271
1100 271
1100 256
1082 256
4 8 15 0 0 0 0 22 20 0 0 4
1143 256
1081 256
1081 256
1082 256
3 7 13 0 0 0 0 22 20 0 0 4
1143 247
1081 247
1081 247
1082 247
2 6 14 0 0 0 0 22 20 0 0 4
1143 238
1081 238
1081 238
1082 238
5 1 16 0 0 4224 0 20 22 0 0 2
1082 229
1143 229
1 3 17 0 0 4224 0 4 3 0 0 2
165 615
118 615
0 3 18 0 0 4096 0 0 26 30 0 5
405 361
405 524
262 524
262 567
281 567
3 3 19 0 0 16512 0 16 8 0 0 6
1476 434
1480 434
1480 433
1484 433
1484 249
1527 249
0 3 20 0 0 4224 0 0 20 42 0 4
1269 349
999 349
999 247
1012 247
0 3 18 0 0 4224 0 0 36 71 0 4
702 361
358 361
358 265
381 265
2 2 21 0 0 4224 0 4 5 0 0 2
201 615
213 615
3 4 22 0 0 8320 0 5 26 0 0 4
258 606
262 606
262 576
287 576
0 1 6 0 0 4224 0 0 5 99 0 4
287 451
82 451
82 597
213 597
0 2 23 0 0 12416 0 0 3 100 0 5
227 415
227 416
22 416
22 624
72 624
5 1 24 0 0 4224 0 26 2 0 0 2
311 606
311 625
3 2 25 0 0 4224 0 25 26 0 0 2
260 558
287 558
0 3 26 0 0 8192 0 0 12 38 0 3
1533 234
1510 234
1510 314
1 2 26 0 0 0 0 8 8 0 0 2
1533 231
1533 240
1 1 27 0 0 12416 0 37 16 0 0 4
1402 436
1411 436
1411 434
1428 434
2 0 28 0 0 12416 0 13 0 0 48 4
1274 398
1274 402
1353 402
1353 249
0 1 29 0 0 4224 0 0 13 47 0 4
1348 258
1348 417
1256 417
1256 398
3 0 20 0 0 0 0 13 0 0 43 5
1265 353
1265 349
1269 349
1269 245
1278 245
1 2 20 0 0 0 0 9 9 0 0 2
1278 240
1278 249
4 0 30 0 0 12416 0 9 0 0 46 5
1272 267
1263 267
1263 282
1344 282
1344 267
3 0 26 0 0 12416 0 9 0 0 37 6
1272 258
1252 258
1252 335
1453 335
1453 278
1510 278
4 8 30 0 0 0 0 11 9 0 0 2
1362 267
1342 267
3 7 29 0 0 0 0 11 9 0 0 2
1362 258
1342 258
2 6 28 0 0 0 0 11 9 0 0 2
1362 249
1342 249
1 5 31 0 0 4224 0 11 9 0 0 2
1362 240
1342 240
0 1 32 0 0 8320 0 0 12 56 0 4
1635 249
1635 377
1501 377
1501 359
0 2 33 0 0 4224 0 0 12 54 0 4
1625 231
1625 367
1519 367
1519 359
7 7 34 0 0 4224 0 6 7 0 0 3
1709 231
1744 231
1744 197
0 4 35 0 0 8320 0 0 8 57 0 4
1608 258
1608 302
1527 302
1527 258
1 5 33 0 0 0 0 6 8 0 0 2
1639 231
1597 231
2 6 36 0 0 4224 0 6 8 0 0 2
1639 240
1597 240
3 7 32 0 0 0 0 6 8 0 0 2
1639 249
1597 249
4 8 35 0 0 0 0 6 8 0 0 2
1639 258
1597 258
7 7 37 0 0 8320 0 11 10 0 0 3
1432 240
1477 240
1477 194
8 6 38 0 0 8320 0 11 10 0 0 3
1432 249
1471 249
1471 194
9 5 39 0 0 8320 0 11 10 0 0 3
1432 258
1465 258
1465 194
10 4 40 0 0 8320 0 11 10 0 0 3
1432 267
1459 267
1459 194
11 3 41 0 0 8320 0 11 10 0 0 3
1432 276
1453 276
1453 194
12 2 42 0 0 8320 0 11 10 0 0 3
1432 285
1447 285
1447 194
13 1 43 0 0 8320 0 11 10 0 0 3
1432 294
1441 294
1441 194
8 6 44 0 0 8320 0 6 7 0 0 3
1709 240
1738 240
1738 197
9 5 45 0 0 8320 0 6 7 0 0 3
1709 249
1732 249
1732 197
10 4 46 0 0 8320 0 6 7 0 0 3
1709 258
1726 258
1726 197
11 3 47 0 0 8320 0 6 7 0 0 3
1709 267
1720 267
1720 197
12 2 48 0 0 12416 0 6 7 0 0 4
1709 276
1709 277
1714 277
1714 197
13 1 49 0 0 8320 0 6 7 0 0 3
1709 285
1708 285
1708 197
3 0 18 0 0 0 0 14 0 0 72 2
702 361
702 240
1 2 18 0 0 0 0 19 19 0 0 7
728 247
728 240
702 240
702 240
715 240
715 256
728 256
3 7 10 0 0 0 0 17 19 0 0 2
858 265
792 265
2 6 11 0 0 0 0 17 19 0 0 2
858 256
792 256
1 5 50 0 0 4224 0 17 19 0 0 2
858 247
792 247
7 7 51 0 0 4224 0 22 21 0 0 3
1213 229
1257 229
1257 203
7 7 52 0 0 4224 0 17 18 0 0 3
928 247
976 247
976 209
8 6 53 0 0 8320 0 17 18 0 0 3
928 256
970 256
970 209
9 5 54 0 0 8320 0 17 18 0 0 3
928 265
964 265
964 209
10 4 55 0 0 8320 0 17 18 0 0 3
928 274
958 274
958 209
11 3 56 0 0 8320 0 17 18 0 0 3
928 283
952 283
952 209
12 2 57 0 0 8320 0 17 18 0 0 3
928 292
946 292
946 209
13 1 58 0 0 8320 0 17 18 0 0 3
928 301
940 301
940 209
8 6 59 0 0 4224 0 22 21 0 0 3
1213 238
1251 238
1251 203
9 5 60 0 0 8320 0 22 21 0 0 3
1213 247
1245 247
1245 203
10 4 61 0 0 8320 0 22 21 0 0 3
1213 256
1239 256
1239 203
11 3 62 0 0 8320 0 22 21 0 0 3
1213 265
1233 265
1233 203
12 2 63 0 0 8320 0 22 21 0 0 3
1213 274
1227 274
1227 203
13 1 64 0 0 8320 0 22 21 0 0 3
1213 283
1221 283
1221 203
0 2 5 0 0 0 0 0 25 101 0 5
207 273
207 429
104 429
104 567
215 567
0 1 7 0 0 8320 0 0 23 8 0 5
354 439
354 438
93 438
93 524
151 524
3 1 65 0 0 8320 0 23 25 0 0 4
196 533
199 533
199 549
215 549
1 7 66 0 0 8320 0 24 26 0 0 3
551 550
551 558
335 558
0 3 67 0 0 4224 0 0 30 95 0 4
345 355
141 355
141 249
147 249
3 2 67 0 0 0 0 33 27 0 0 2
345 369
345 336
3 1 68 0 0 8192 0 29 27 0 0 4
278 366
278 342
327 342
327 336
0 0 68 0 0 4224 0 0 0 96 102 4
278 342
94 342
94 235
153 235
2 3 69 0 0 8320 0 36 27 0 0 4
387 256
387 253
336 253
336 290
2 3 6 0 0 0 0 29 28 0 0 3
287 411
287 470
323 470
1 0 23 0 0 0 0 29 0 0 104 4
269 411
269 415
227 415
227 249
0 4 5 0 0 0 0 0 30 103 0 5
223 258
223 273
145 273
145 258
147 258
2 1 68 0 0 0 0 30 30 0 0 6
153 240
153 235
155 235
155 235
153 235
153 231
4 8 5 0 0 0 0 31 30 0 0 2
230 258
217 258
3 7 23 0 0 0 0 31 30 0 0 2
230 249
217 249
2 6 70 0 0 4224 0 31 30 0 0 2
230 240
217 240
1 5 71 0 0 4224 0 31 30 0 0 2
230 231
217 231
7 7 72 0 0 4224 0 31 32 0 0 3
300 231
338 231
338 219
8 6 73 0 0 4224 0 31 32 0 0 3
300 240
332 240
332 219
9 5 74 0 0 8320 0 31 32 0 0 3
300 249
326 249
326 219
10 4 75 0 0 8320 0 31 32 0 0 3
300 258
320 258
320 219
11 3 76 0 0 8320 0 31 32 0 0 3
300 267
314 267
314 219
12 2 77 0 0 8320 0 31 32 0 0 3
300 276
308 276
308 219
13 1 78 0 0 8320 0 31 32 0 0 3
300 285
302 285
302 219
2 1 69 0 0 0 0 36 36 0 0 2
387 256
387 247
7 3 7 0 0 0 0 36 34 0 0 2
451 265
492 265
7 7 79 0 0 4224 0 34 35 0 0 3
562 247
596 247
596 215
8 6 80 0 0 8320 0 34 35 0 0 3
562 256
590 256
590 215
9 5 81 0 0 8320 0 34 35 0 0 3
562 265
584 265
584 215
10 4 82 0 0 8320 0 34 35 0 0 3
562 274
578 274
578 215
11 3 83 0 0 8320 0 34 35 0 0 3
562 283
572 283
572 215
12 2 84 0 0 8320 0 34 35 0 0 3
562 292
566 292
566 215
13 1 85 0 0 8320 0 34 35 0 0 3
562 301
560 301
560 215
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
